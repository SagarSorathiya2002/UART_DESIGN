package transaction;

class transaction;
  
  rand logic [7:0] tx_byte;
       logic [7:0] rx_byte;
       logic [1:0] baud_sel;
       logic tx_enable;
       logic rx_bussy,rx_error,rx_valid;
       logic TX_VALID,TX_BUSSY;
       logic rst; 
       
  
endclass 
endpackage 