package file;

`include"transaction.sv"
`include"UART_driver.sv"
`include"UART_generator.sv"
`include"UART_monitor.sv"

endpackage
